// Registers for elevator floors
module register( );

endmodule //register
